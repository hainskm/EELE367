entity add_n_sub_8bit is
	port (A, B : in std_logic_vector(7 downto 0);
	      ADDn_SUB : in std_logic;
	      Sum_DIFF : out std_logic_vector(7 downto 0);
	      Cout_Bout : out std_logic;
	      Vout : out std_logic);
end entity;

architecture add_n_sub_8bit_arch of add_n_sub_8bit is

	begin

end architecture;
