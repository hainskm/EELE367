library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity fsm2_behavioral is
	port (Clock, Reset : in std_logic;
	      Din	   : in std_logic;
	      Dout	   : out std_logic);
end entity;

architecture fsm2_behavioral_arch of fsm2_behavioral is
	type State_Type is (S0, S1, S2, S3);
	signal curr_state, next_state : State_Type;

	begin
		STATE_MEMORY : process (Clock, Reset)
			begin
				if (Reset = '0') then
					curr_state <= S0;
				elsif (Clock'event and Clock = '1') then
					curr_state <= next_state;
				end if;
		end process;
	
		NEXT_STATE_LOGIC : process(curr_state, Din)
			begin
				case (curr_state) is
					when S0 => if (Din = '1') then	
							next_state <= S1;
						   else
							next_state <= S0;
						   end if;
					when S1 => if (Din = '1') then	
							next_state <= S3;
						   else
							next_state <= S2;
						   end if;
					when s2 => if (Din = '1') then	
							next_state <= S3;
						   else
							next_state <= S0;
						   end if;
					when s3 => if (Din = '1') then	
							next_state <= S0;
						   else
							next_state <= S3;
						   end if;
				end case;
		end process;

		OUTPUT_LOGIC : process(curr_state, Din)
			begin
				case(curr_state) is
					when S0 => if (Din = '1') then	
							Dout <= '1';
						   else
							Dout <= '0';
						   end if;
					when S1 => if (Din = '1') then	
							Dout <= '0';
						   else
							Dout <= '1';
						   end if;
					when S2 => if (Din = '1') then	
							Dout <= '1';
						   else
							Dout <= '0';
						   end if;
					when S3 => if (Din = '1') then	
							Dout <= '1';
						   else
							Dout <= '0';
						   end if;
				end case;
		end process;
end architecture;
